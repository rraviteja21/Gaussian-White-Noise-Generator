
`include "def.v"

module ln_mul( x_e,			// input to log function
	       y_e );			// output of log function

input [48 : 0]x_e;
output [31:0]y_e;		
wire [7:0]x_e_a;
wire [48 : 0]x_e_b;		

wire [12 : 0] C2;			// coefficients of piecewise polynomial.
wire [21: 0]  C1;
wire [29:0]   C0;

assign x_e_a = x_e[48:41];				// range reduction
assign x_e_b = x_e[40:0] << 8;			

ln_poly ln_poly0(.x_e_a(x_e_a),
				 .C2_ret(C2),
				 .C1_ret(C1),
				 .C0_ret(C0) );
				 
/*Multiplies the coefficients with the input and produces the output*/
myMultiplier_ln2 myMultiplier_ln2_0(  .x(x_e_b),				
									  .C2(C2),
									  .C1(C1),
									  .C0(C0),
									  .result(y_e));	
endmodule


/******************************* This module acts as the look up for the logarithm and outputs the required coefficients*****************************/

module ln_poly( x_e_a,
		        C2_ret,
		        C1_ret,
		        C0_ret);
input [7:0]x_e_a;
output [12 : 0]        C2_ret;
output [21: 0]        C1_ret;
output [29:0]        C0_ret;

reg [12 : 0] C2;
reg [21: 0]  C1;
reg [29:0]   C0;


assign C2_ret = C2;
assign C1_ret = C1;
assign C0_ret = C0;

always @(*)
begin
	case(x_e_a)
		
8'd0:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111111111000000
;
      C0 <= 30'b101000000001111111110001010111
;
     end
8'd1:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111111100000010
;
      C0 <= 30'b101000001101111011010011001101
;
     end
8'd2:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111111001000110
;
      C0 <= 30'b101000011001110000111011011110
;
     end
8'd3:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111110110001011
;
      C0 <= 30'b101000100101100000101111000000
;
     end
8'd4:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111110011010011
;
      C0 <= 30'b101000110001001010110010100010
;
     end
8'd5:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111110000011100
;
      C0 <= 30'b101000111100101111001010110001
;
     end
8'd6:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111101101100111
;
      C0 <= 30'b101001001000001101111100010010
;
     end
8'd7:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111101010110101
;
      C0 <= 30'b101001010011100111001011100111
;
     end
8'd8:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111101000000011
;
      C0 <= 30'b101001011110111010111101001100
;
     end
8'd9:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111100101010100
;
      C0 <= 30'b101001101010001001010101011001
;
     end
8'd10:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111100010100110
;
      C0 <= 30'b101001110101010010011000100000
;
     end
8'd11:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111011111111011
;
      C0 <= 30'b101010000000010110001010110000
;
     end
8'd12:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111011101010000
;
      C0 <= 30'b101010001011010100110000010010
;
     end
8'd13:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111011010101000
;
      C0 <= 30'b101010010110001110001101001011
;
     end
8'd14:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111011000000001
;
      C0 <= 30'b101010100001000010100101011101
;
     end
8'd15:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111010101011100
;
      C0 <= 30'b101010101011110001111101000100
;
     end
8'd16:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111010010111000
;
      C0 <= 30'b101010110110011100010111111001
;
     end
8'd17:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111010000010110
;
      C0 <= 30'b101011000001000001111001110001
;
     end
8'd18:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111001101110110
;
      C0 <= 30'b101011001011100010100110011011
;
     end
8'd19:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111001011010111
;
      C0 <= 30'b101011010101111110100001100101
;
     end
8'd20:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111001000111001
;
      C0 <= 30'b101011100000010101101110110111
;
     end
8'd21:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111000110011101
;
      C0 <= 30'b101011101010101000010001110110
;
     end
8'd22:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111000100000011
;
      C0 <= 30'b101011110100110110001110000101
;
     end
8'd23:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000111000001101010
;
      C0 <= 30'b101011111110111111100110111111
;
     end
8'd24:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110111111010011
;
      C0 <= 30'b101100001001000100100000000001
;
     end
8'd25:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110111100111100
;
      C0 <= 30'b101100010011000100111100100000
;
     end
8'd26:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110111010101000
;
      C0 <= 30'b101100011101000000111111110001
;
     end
8'd27:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110111000010100
;
      C0 <= 30'b101100100110111000101101000010
;
     end
8'd28:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110110110000011
;
      C0 <= 30'b101100110000101100000111100010
;
     end
8'd29:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110110011110010
;
      C0 <= 30'b101100111010011011010010011001
;
     end
8'd30:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110110001100011
;
      C0 <= 30'b101101000100000110010000101111
;
     end
8'd31:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110101111010101
;
      C0 <= 30'b101101001101101101000101100110
;
     end
8'd32:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110101101001000
;
      C0 <= 30'b101101010111001111110100000000
;
     end
8'd33:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110101010111101
;
      C0 <= 30'b101101100000101110011110111001
;
     end
8'd34:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110101000110011
;
      C0 <= 30'b101101101010001001001001001101
;
     end
8'd35:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110100110101010
;
      C0 <= 30'b101101110011011111110101110010
;
     end
8'd36:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110100100100010
;
      C0 <= 30'b101101111100110010100111011111
;
     end
8'd37:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110100010011100
;
      C0 <= 30'b101110000110000001100001000100
;
     end
8'd38:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110100000010111
;
      C0 <= 30'b101110001111001100100101010011
;
     end
8'd39:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110011110010011
;
      C0 <= 30'b101110011000010011110110110111
;
     end
8'd40:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110011100010000
;
      C0 <= 30'b101110100001010111011000011011
;
     end
8'd41:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110011010001110
;
      C0 <= 30'b101110101010010111001100100111
;
     end
8'd42:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110011000001101
;
      C0 <= 30'b101110110011010011010110000000
;
     end
8'd43:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110010110001110
;
      C0 <= 30'b101110111100001011110111001001
;
     end
8'd44:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110010100010000
;
      C0 <= 30'b101111000101000000110010100011
;
     end
8'd45:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110010010010011
;
      C0 <= 30'b101111001101110010001010101011
;
     end
8'd46:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110010000010110
;
      C0 <= 30'b101111010110100000000001111101
;
     end
8'd47:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110001110011011
;
      C0 <= 30'b101111011111001010011010110011
;
     end
8'd48:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110001100100001
;
      C0 <= 30'b101111100111110001010111100100
;
     end
8'd49:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110001010101001
;
      C0 <= 30'b101111110000010100111010100110
;
     end
8'd50:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110001000110001
;
      C0 <= 30'b101111111000110101000110001011
;
     end
8'd51:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110000110111010
;
      C0 <= 30'b110000000001010001111100100100
;
     end
8'd52:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110000101000100
;
      C0 <= 30'b110000001001101011011111111111
;
     end
8'd53:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110000011001111
;
      C0 <= 30'b110000010010000001110010101011
;
     end
8'd54:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000110000001011011
;
      C0 <= 30'b110000011010010100110110110001
;
     end
8'd55:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101111111101000
;
      C0 <= 30'b110000100010100100101110011010
;
     end
8'd56:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101111101110110
;
      C0 <= 30'b110000101010110001011011101100
;
     end
8'd57:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101111100000101
;
      C0 <= 30'b110000110010111011000000101110
;
     end
8'd58:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101111010010101
;
      C0 <= 30'b110000111011000001011111100010
;
     end
8'd59:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101111000100110
;
      C0 <= 30'b110001000011000100111010001010
;
     end
8'd60:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101110110111000
;
      C0 <= 30'b110001001011000101010010100100
;
     end
8'd61:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101110101001011
;
      C0 <= 30'b110001010011000010101010101111
;
     end
8'd62:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101110011011110
;
      C0 <= 30'b110001011010111101000100100110
;
     end
8'd63:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101110001110011
;
      C0 <= 30'b110001100010110100100010000100
;
     end
8'd64:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101110000001000
;
      C0 <= 30'b110001101010101001000101000001
;
     end
8'd65:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101101110011110
;
      C0 <= 30'b110001110010011010101111010101
;
     end
8'd66:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101101100110110
;
      C0 <= 30'b110001111010001001100010110100
;
     end
8'd67:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101101011001110
;
      C0 <= 30'b110010000001110101100001010011
;
     end
8'd68:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101101001100110
;
      C0 <= 30'b110010001001011110101100100011
;
     end
8'd69:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101101000000000
;
      C0 <= 30'b110010010001000101000110010110
;
     end
8'd70:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101100110011010
;
      C0 <= 30'b110010011000101000110000011001
;
     end
8'd71:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101100100110110
;
      C0 <= 30'b110010100000001001101100011100
;
     end
8'd72:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101100011010010
;
      C0 <= 30'b110010100111100111111100001010
;
     end
8'd73:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101100001101110
;
      C0 <= 30'b110010101111000011100001001110
;
     end
8'd74:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101100000001100
;
      C0 <= 30'b110010110110011100011101010001
;
     end
8'd75:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101011110101010
;
      C0 <= 30'b110010111101110010110001111010
;
     end
8'd76:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101011101001010
;
      C0 <= 30'b110011000101000110100000110010
;
     end
8'd77:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101011011101010
;
      C0 <= 30'b110011001100010111101011011101
;
     end
8'd78:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101011010001010
;
      C0 <= 30'b110011010011100110010011011110
;
     end
8'd79:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101011000101100
;
      C0 <= 30'b110011011010110010011010011001
;
     end
8'd80:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010111001110
;
      C0 <= 30'b110011100001111100000001101110
;
     end
8'd81:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010101110001
;
      C0 <= 30'b110011101001000011001010111111
;
     end
8'd82:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010100010100
;
      C0 <= 30'b110011110000000111110111101000
;
     end
8'd83:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010010111000
;
      C0 <= 30'b110011110111001010001001001001
;
     end
8'd84:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010001011101
;
      C0 <= 30'b110011111110001010000000111110
;
     end
8'd85:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101010000000011
;
      C0 <= 30'b110100000101000111100000100001
;
     end
8'd86:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101001110101001
;
      C0 <= 30'b110100001100000010101001001101
;
     end
8'd87:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101001101010000
;
      C0 <= 30'b110100010010111011011100011011
;
     end
8'd88:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101001011111000
;
      C0 <= 30'b110100011001110001111011100011
;
     end
8'd89:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101001010100000
;
      C0 <= 30'b110100100000100110000111111011
;
     end
8'd90:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101001001001001
;
      C0 <= 30'b110100100111011000000010111000
;
     end
8'd91:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000111110011
;
      C0 <= 30'b110100101110000111101101110000
;
     end
8'd92:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000110011101
;
      C0 <= 30'b110100110100110101001001110110
;
     end
8'd93:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000101001000
;
      C0 <= 30'b110100111011100000011000011101
;
     end
8'd94:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000011110100
;
      C0 <= 30'b110101000010001001011010110101
;
     end
8'd95:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000010100000
;
      C0 <= 30'b110101001000110000010010001111
;
     end
8'd96:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000101000001001101
;
      C0 <= 30'b110101001111010100111111111010
;
     end
8'd97:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111111111010
;
      C0 <= 30'b110101010101110111100101000110
;
     end
8'd98:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111110101000
;
      C0 <= 30'b110101011100011000000010111111
;
     end
8'd99:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111101010111
;
      C0 <= 30'b110101100010110110011010110001
;
     end
8'd100:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111100000110
;
      C0 <= 30'b110101101001010010101101101010
;
     end
8'd101:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111010110110
;
      C0 <= 30'b110101101111101100111100110011
;
     end
8'd102:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111001100110
;
      C0 <= 30'b110101110110000101001001010110
;
     end
8'd103:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100111000010111
;
      C0 <= 30'b110101111100011011010100011011
;
     end
8'd104:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110111001001
;
      C0 <= 30'b110110000010101111011111001100
;
     end
8'd105:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110101111011
;
      C0 <= 30'b110110001001000001101010101111
;
     end
8'd106:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110100101110
;
      C0 <= 30'b110110001111010001111000001010
;
     end
8'd107:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110011100001
;
      C0 <= 30'b110110010101100000001000100011
;
     end
8'd108:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110010010101
;
      C0 <= 30'b110110011011101100011100111111
;
     end
8'd109:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100110001001001
;
      C0 <= 30'b110110100001110110110110100001
;
     end
8'd110:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101111111110
;
      C0 <= 30'b110110100111111111010110001100
;
     end
8'd111:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101110110011
;
      C0 <= 30'b110110101110000101111101000011
;
     end
8'd112:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101101101001
;
      C0 <= 30'b110110110100001010101100000111
;
     end
8'd113:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101100011111
;
      C0 <= 30'b110110111010001101100100011001
;
     end
8'd114:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101011010110
;
      C0 <= 30'b110111000000001110100110111001
;
     end
8'd115:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101010001101
;
      C0 <= 30'b110111000110001101110100100110
;
     end
8'd116:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100101001000101
;
      C0 <= 30'b110111001100001011001110011110
;
     end
8'd117:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100111111110
;
      C0 <= 30'b110111010010000110110101011111
;
     end
8'd118:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100110110111
;
      C0 <= 30'b110111011000000000101010100110
;
     end
8'd119:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100101110000
;
      C0 <= 30'b110111011101111000101110110000
;
     end
8'd120:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100100101010
;
      C0 <= 30'b110111100011101111000010111001
;
     end
8'd121:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100011100100
;
      C0 <= 30'b110111101001100011100111111010
;
     end
8'd122:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100010011111
;
      C0 <= 30'b110111101111010110011110101111
;
     end
8'd123:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100001011010
;
      C0 <= 30'b110111110101000111101000010001
;
     end
8'd124:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100100000010110
;
      C0 <= 30'b110111111010110111000101011001
;
     end
8'd125:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011111010010
;
      C0 <= 30'b111000000000100100110111000000
;
     end
8'd126:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011110001111
;
      C0 <= 30'b111000000110010000111101111101
;
     end
8'd127:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011101001100
;
      C0 <= 30'b111000001011111011011011000111
;
     end
8'd128:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011100001010
;
      C0 <= 30'b111000010001100100001111010101
;
     end
8'd129:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011011001000
;
      C0 <= 30'b111000010111001011011011011100
;
     end
8'd130:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011010000110
;
      C0 <= 30'b111000011100110001000000010011
;
     end
8'd131:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011001000101
;
      C0 <= 30'b111000100010010100111110101100
;
     end
8'd132:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100011000000100
;
      C0 <= 30'b111000100111110111010111011110
;
     end
8'd133:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010111000100
;
      C0 <= 30'b111000101101011000001011011011
;
     end
8'd134:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010110000100
;
      C0 <= 30'b111000110010110111011011010101
;
     end
8'd135:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010101000101
;
      C0 <= 30'b111000111000010101001000000001
;
     end
8'd136:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010100000110
;
      C0 <= 30'b111000111101110001010010001110
;
     end
8'd137:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010011000111
;
      C0 <= 30'b111001000011001011111010110000
;
     end
8'd138:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010010001001
;
      C0 <= 30'b111001001000100101000010010110
;
     end
8'd139:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010001001011
;
      C0 <= 30'b111001001101111100101001110000
;
     end
8'd140:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100010000001110
;
      C0 <= 30'b111001010011010010110001101111
;
     end
8'd141:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001111010001
;
      C0 <= 30'b111001011000100111011011000001
;
     end
8'd142:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001110010100
;
      C0 <= 30'b111001011101111010100110010110
;
     end
8'd143:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001101011000
;
      C0 <= 30'b111001100011001100010100011100
;
     end
8'd144:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001100011100
;
      C0 <= 30'b111001101000011100100101111111
;
     end
8'd145:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001011100000
;
      C0 <= 30'b111001101101101011011011101110
;
     end
8'd146:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001010100101
;
      C0 <= 30'b111001110010111000110110010110
;
     end
8'd147:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001001101011
;
      C0 <= 30'b111001111000000100110110100001
;
     end
8'd148:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100001000110000
;
      C0 <= 30'b111001111101001111011100111101
;
     end
8'd149:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000111110110
;
      C0 <= 30'b111010000010011000101010010101
;
     end
8'd150:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000110111101
;
      C0 <= 30'b111010000111100000011111010011
;
     end
8'd151:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000110000100
;
      C0 <= 30'b111010001100100110111100100010
;
     end
8'd152:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000101001011
;
      C0 <= 30'b111010010001101100000010101100
;
     end
8'd153:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000100010010
;
      C0 <= 30'b111010010110101111110010011011
;
     end
8'd154:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000011011010
;
      C0 <= 30'b111010011011110010001100010111
;
     end
8'd155:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000010100010
;
      C0 <= 30'b111010100000110011010001001001
;
     end
8'd156:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000001101011
;
      C0 <= 30'b111010100101110011000001011010
;
     end
8'd157:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000100000000110100
;
      C0 <= 30'b111010101010110001011101110010
;
     end
8'd158:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111111111101
;
      C0 <= 30'b111010101111101110100110110111
;
     end
8'd159:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111111000110
;
      C0 <= 30'b111010110100101010011101010010
;
     end
8'd160:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111110010000
;
      C0 <= 30'b111010111001100101000001101000
;
     end
8'd161:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111101011010
;
      C0 <= 30'b111010111110011110010100100000
;
     end
8'd162:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111100100101
;
      C0 <= 30'b111011000011010110010110100000
;
     end
8'd163:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111011110000
;
      C0 <= 30'b111011001000001101001000001101
;
     end
8'd164:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111010111011
;
      C0 <= 30'b111011001101000010101010001101
;
     end
8'd165:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111010000110
;
      C0 <= 30'b111011010001110110111101000011
;
     end
8'd166:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111001010010
;
      C0 <= 30'b111011010110101010000001010110
;
     end
8'd167:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011111000011110
;
      C0 <= 30'b111011011011011011110111100111
;
     end
8'd168:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110111101011
;
      C0 <= 30'b111011100000001100100000011100
;
     end
8'd169:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110110111000
;
      C0 <= 30'b111011100100111011111100011000
;
     end
8'd170:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110110000101
;
      C0 <= 30'b111011101001101010001011111101
;
     end
8'd171:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110101010010
;
      C0 <= 30'b111011101110010111001111101101
;
     end
8'd172:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110100100000
;
      C0 <= 30'b111011110011000011001000001100
;
     end
8'd173:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110011101110
;
      C0 <= 30'b111011110111101101110101111011
;
     end
8'd174:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110010111100
;
      C0 <= 30'b111011111100010111011001011100
;
     end
8'd175:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110010001010
;
      C0 <= 30'b111100000000111111110011010000
;
     end
8'd176:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110001011001
;
      C0 <= 30'b111100000101100111000011111000
;
     end
8'd177:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011110000101000
;
      C0 <= 30'b111100001010001101001011110101
;
     end
8'd178:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101111111000
;
      C0 <= 30'b111100001110110010001011100110
;
     end
8'd179:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101111000111
;
      C0 <= 30'b111100010011010110000011101100
;
     end
8'd180:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101110010111
;
      C0 <= 30'b111100010111111000110100100110
;
     end
8'd181:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101101101000
;
      C0 <= 30'b111100011100011010011110110100
;
     end
8'd182:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101100111000
;
      C0 <= 30'b111100100000111011000010110110
;
     end
8'd183:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101100001001
;
      C0 <= 30'b111100100101011010100001001000
;
     end
8'd184:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101011011010
;
      C0 <= 30'b111100101001111000111010001011
;
     end
8'd185:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101010101011
;
      C0 <= 30'b111100101110010110001110011101
;
     end
8'd186:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101001111101
;
      C0 <= 30'b111100110010110010011110011010
;
     end
8'd187:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101001001111
;
      C0 <= 30'b111100110111001101101010100001
;
     end
8'd188:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011101000100001
;
      C0 <= 30'b111100111011100111110011010000
;
     end
8'd189:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100111110011
;
      C0 <= 30'b111101000000000000111001000010
;
     end
8'd190:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100111000110
;
      C0 <= 30'b111101000100011000111100010101
;
     end
8'd191:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100110011001
;
      C0 <= 30'b111101001000101111111101100110
;
     end
8'd192:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100101101100
;
      C0 <= 30'b111101001101000101111101010001
;
     end
8'd193:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100101000000
;
      C0 <= 30'b111101010001011010111011110001
;
     end
8'd194:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100100010011
;
      C0 <= 30'b111101010101101110111001100010
;
     end
8'd195:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100011100111
;
      C0 <= 30'b111101011010000001110111000001
;
     end
8'd196:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100010111011
;
      C0 <= 30'b111101011110010011110100100111
;
     end
8'd197:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100010010000
;
      C0 <= 30'b111101100010100100110010110000
;
     end
8'd198:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100001100100
;
      C0 <= 30'b111101100110110100110001110111
;
     end
8'd199:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100000111001
;
      C0 <= 30'b111101101011000011110010010110
;
     end
8'd200:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011100000001111
;
      C0 <= 30'b111101101111010001110100100111
;
     end
8'd201:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011111100100
;
      C0 <= 30'b111101110011011110111001000101
;
     end
8'd202:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011110111010
;
      C0 <= 30'b111101110111101011000000001000
;
     end
8'd203:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011110001111
;
      C0 <= 30'b111101111011110110001010001011
;
     end
8'd204:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011101100101
;
      C0 <= 30'b111110000000000000010111100111
;
     end
8'd205:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011100111100
;
      C0 <= 30'b111110000100001001101000110100
;
     end
8'd206:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011100010010
;
      C0 <= 30'b111110001000010001111110001100
;
     end
8'd207:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011011101001
;
      C0 <= 30'b111110001100011001011000001000
;
     end
8'd208:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011011000000
;
      C0 <= 30'b111110010000011111110110111110
;
     end
8'd209:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011010010111
;
      C0 <= 30'b111110010100100101011011001001
;
     end
8'd210:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011001101111
;
      C0 <= 30'b111110011000101010000100111111
;
     end
8'd211:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011001000110
;
      C0 <= 30'b111110011100101101110100111000
;
     end
8'd212:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011011000011110
;
      C0 <= 30'b111110100000110000101011001100
;
     end
8'd213:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010111110110
;
      C0 <= 30'b111110100100110010101000010010
;
     end
8'd214:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010111001110
;
      C0 <= 30'b111110101000110011101100100010
;
     end
8'd215:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010110100111
;
      C0 <= 30'b111110101100110011111000010001
;
     end
8'd216:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010110000000
;
      C0 <= 30'b111110110000110011001011110111
;
     end
8'd217:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010101011001
;
      C0 <= 30'b111110110100110001100111101011
;
     end
8'd218:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010100110010
;
      C0 <= 30'b111110111000101111001100000001
;
     end
8'd219:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010100001011
;
      C0 <= 30'b111110111100101011111001010010
;
     end
8'd220:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010011100101
;
      C0 <= 30'b111111000000100111101111110010
;
     end
8'd221:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010010111110
;
      C0 <= 30'b111111000100100010101111110111
;
     end
8'd222:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010010011000
;
      C0 <= 30'b111111001000011100111001110110
;
     end
8'd223:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010001110010
;
      C0 <= 30'b111111001100010110001110000110
;
     end
8'd224:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010001001101
;
      C0 <= 30'b111111010000001110101100111011
;
     end
8'd225:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010000100111
;
      C0 <= 30'b111111010100000110010110101010
;
     end
8'd226:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011010000000010
;
      C0 <= 30'b111111010111111101001011100111
;
     end
8'd227:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001111011101
;
      C0 <= 30'b111111011011110011001100001000
;
     end
8'd228:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001110111000
;
      C0 <= 30'b111111011111101000011000100001
;
     end
8'd229:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001110010011
;
      C0 <= 30'b111111100011011100110001000111
;
     end
8'd230:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001101101111
;
      C0 <= 30'b111111100111010000010110001100
;
     end
8'd231:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001101001011
;
      C0 <= 30'b111111101011000011001000000101
;
     end
8'd232:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001100100110
;
      C0 <= 30'b111111101110110101000111000110
;
     end
8'd233:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001100000011
;
      C0 <= 30'b111111110010100110010011100011
;
     end
8'd234:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001011011111
;
      C0 <= 30'b111111110110010110101101101110
;
     end
8'd235:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001010111011
;
      C0 <= 30'b111111111010000110010101111011
;
     end
8'd236:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001010011000
;
      C0 <= 30'b111111111101110101001100011110
;
     end
8'd237:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001001110101
;
      C0 <= 30'b000000000001100011010001101000
;
     end
8'd238:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001001010010
;
      C0 <= 30'b000000000101010000100101101101
;
     end
8'd239:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001000101111
;
      C0 <= 30'b000000001000111101001000111111
;
     end
8'd240:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011001000001100
;
      C0 <= 30'b000000001100101000111011110010
;
     end
8'd241:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000111101001
;
      C0 <= 30'b000000010000010011111110010110
;
     end
8'd242:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000111000111
;
      C0 <= 30'b000000010011111110010000111110
;
     end
8'd243:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000110100101
;
      C0 <= 30'b000000010111100111110011111101
;
     end
8'd244:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000110000011
;
      C0 <= 30'b000000011011010000100111100011
;
     end
8'd245:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000101100001
;
      C0 <= 30'b000000011110111000101100000011
;
     end
8'd246:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000101000000
;
      C0 <= 30'b000000100010100000000001101111
;
     end
8'd247:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000100011110
;
      C0 <= 30'b000000100110000110101000110111
;
     end
8'd248:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000011111101
;
      C0 <= 30'b000000101001101100100001101101
;
     end
8'd249:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000011011100
;
      C0 <= 30'b000000101101010001101100100001
;
     end
8'd250:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000010111011
;
      C0 <= 30'b000000110000110110001001100110
;
     end
8'd251:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000010011010
;
      C0 <= 30'b000000110100011001111001001100
;
     end
8'd252:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000001111001
;
      C0 <= 30'b000000110111111100111011100011
;
     end
8'd253:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000001011001
;
      C0 <= 30'b000000111011011111010000111100
;
     end
8'd254:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000000111000
;
      C0 <= 30'b000000111111000000111001101000
;
     end
8'd255:
      begin
      C2 <= 13'b0000000000000
;
      C1 <= 22'b0000000011000000011000
;
      C0 <= 30'b000001000010100001110101110110
;
     end
 

	default:
	begin				// default case
		C2 <= 13'b0;
		C1 <= 22'b0;
		C0 <= 30'b0;
	end
	
 endcase
 end
 endmodule

