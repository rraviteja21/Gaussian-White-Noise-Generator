


module cos_mul( x_g_a,
				x_g_b,
				y_g_a,
				y_g_b);
input [13:0]x_g_a, x_g_b;
output [15:0]y_g_a, y_g_b;

wire [11:0]C1_a;
wire [18:0]C0_a;						   	// coefficients of piecewise polynomial for cos function
wire [11:0]C1_b;
wire [18:0]C0_b;								// coefficients of piecewise polynomial for sin function

																		// gets coefficients for cos function
cos_poly cos_poly_0(.x_g(x_g_a[13:7]),
					.C1_o(C1_a),
					.C0_o(C0_a));
																			// gets coefficients for sin function				
cos_poly sin_poly_1(.x_g(x_g_b[13:7]),
					.C1_o(C1_b),
					.C0_o(C0_b) );

/*Multiplies the coefficients with the input and produces the output*/					
					
myMultiplier_cos myMultiplier_cos( .x_g(x_g_a << 7),
								   .C1(C1_a),
								   .C0(C0_a),
								   .y_g(y_g_a));
								   
myMultiplier_cos myMultiplier_sin( .x_g(x_g_b << 7),
								   .C1(C1_b),
								   .C0(C0_b),
								   .y_g(y_g_b) );
				
endmodule


/******************************* This module acts as the look up for the cos/sine functions and outputs the required coefficients*****************************/
module cos_poly( x_g,
				 C1_o,
				 C0_o);
input [6:0]x_g;				 
output  [11:0]C1_o; // (1,11) signed
output [18:0]C0_o;  // (1,18) unsigned

reg [11:0]C1;
reg [18:0]C0;

assign C1_o = C1;
assign C0_o = C0;

always @(*)
begin
case(x_g)

  7'd0:
     begin
      C1 <= 12'b000000000000
;
      C0 <= 19'b0111111111111111111
;
      end
  7'd1:
     begin
      C1 <= 12'b000000000000
;
      C0 <= 19'b0000000000000000101
;
      end
  7'd2:
     begin
      C1 <= 12'b111111111111
;
      C0 <= 19'b0000000000000111011
;
      end
  7'd3:
     begin
      C1 <= 12'b111111111111
;
      C0 <= 19'b0000000000001100010
;
      end
  7'd4:
     begin
      C1 <= 12'b111111111111
;
      C0 <= 19'b0000000000100111010
;
      end
  7'd5:
     begin
      C1 <= 12'b111111111110
;
      C0 <= 19'b0000000001111000011
;
      end
  7'd6:
     begin
      C1 <= 12'b111111111110
;
      C0 <= 19'b0000000000111111110
;
      end
  7'd7:
     begin
      C1 <= 12'b111111111110
;
      C0 <= 19'b0000000011111101010
;
      end
  7'd8:
     begin
      C1 <= 12'b111111111101
;
      C0 <= 19'b0000000010110001000
;
      end
  7'd9:
     begin
      C1 <= 12'b111111111101
;
      C0 <= 19'b0000000001011011000
;
      end
  7'd10:
     begin
      C1 <= 12'b111111111101
;
      C0 <= 19'b0000000111111011010
;
      end
  7'd11:
     begin
      C1 <= 12'b111111111100
;
      C0 <= 19'b0000000110010001111
;
      end
  7'd12:
     begin
      C1 <= 12'b111111111100
;
      C0 <= 19'b0000000100011110101
;
      end
  7'd13:
     begin
      C1 <= 12'b111111111100
;
      C0 <= 19'b0000000010100001111
;
      end
  7'd14:
     begin
      C1 <= 12'b111111111100
;
      C0 <= 19'b0000000000011011100
;
      end
  7'd15:
     begin
      C1 <= 12'b111111111011
;
      C0 <= 19'b0000001110001011101
;
      end
  7'd16:
     begin
      C1 <= 12'b111111111011
;
      C0 <= 19'b0000001011110010001
;
      end
  7'd17:
     begin
      C1 <= 12'b111111111011
;
      C0 <= 19'b0000001001001111001
;
      end
  7'd18:
     begin
      C1 <= 12'b111111111010
;
      C0 <= 19'b0000000110100010110
;
      end
  7'd19:
     begin
      C1 <= 12'b111111111010
;
      C0 <= 19'b0000000011101101001
;
      end
  7'd20:
     begin
      C1 <= 12'b111111111010
;
      C0 <= 19'b0000000000101110000
;
      end
  7'd21:
     begin
      C1 <= 12'b111111111001
;
      C0 <= 19'b0000011101100101110
;
      end
  7'd22:
     begin
      C1 <= 12'b111111111001
;
      C0 <= 19'b0000011010010100010
;
      end
  7'd23:
     begin
      C1 <= 12'b111111111001
;
      C0 <= 19'b0000010110111001101
;
      end
  7'd24:
     begin
      C1 <= 12'b111111111001
;
      C0 <= 19'b0000010011010101111
;
      end
  7'd25:
     begin
      C1 <= 12'b111111111000
;
      C0 <= 19'b0000001111101001001
;
      end
  7'd26:
     begin
      C1 <= 12'b111111111000
;
      C0 <= 19'b0000001011110011100
;
      end
  7'd27:
     begin
      C1 <= 12'b111111111000
;
      C0 <= 19'b0000000111110101001
;
      end
  7'd28:
     begin
      C1 <= 12'b111111110111
;
      C0 <= 19'b0000000011101101111
;
      end
  7'd29:
     begin
      C1 <= 12'b111111110111
;
      C0 <= 19'b0000111111011101111
;
      end
  7'd30:
     begin
      C1 <= 12'b111111110111
;
      C0 <= 19'b0000111011000101011
;
      end
  7'd31:
     begin
      C1 <= 12'b111111110111
;
      C0 <= 19'b0000110110100100010
;
      end
  7'd32:
     begin
      C1 <= 12'b111111110110
;
      C0 <= 19'b0000110001111010110
;
      end
  7'd33:
     begin
      C1 <= 12'b111111110110
;
      C0 <= 19'b0000101101001001000
;
      end
  7'd34:
     begin
      C1 <= 12'b111111110110
;
      C0 <= 19'b0000101000001110111
;
      end
  7'd35:
     begin
      C1 <= 12'b111111110101
;
      C0 <= 19'b0000100011001100101
;
      end
  7'd36:
     begin
      C1 <= 12'b111111110101
;
      C0 <= 19'b0000011110000010011
;
      end
  7'd37:
     begin
      C1 <= 12'b111111110101
;
      C0 <= 19'b0000011000110000001
;
      end
  7'd38:
     begin
      C1 <= 12'b111111110101
;
      C0 <= 19'b0000010011010110000
;
      end
  7'd39:
     begin
      C1 <= 12'b111111110100
;
      C0 <= 19'b0000001101110100010
;
      end
  7'd40:
     begin
      C1 <= 12'b111111110100
;
      C0 <= 19'b0000001000001010110
;
      end
  7'd41:
     begin
      C1 <= 12'b111111110100
;
      C0 <= 19'b0000000010011001110
;
      end
  7'd42:
     begin
      C1 <= 12'b111111110011
;
      C0 <= 19'b0001111100100001011
;
      end
  7'd43:
     begin
      C1 <= 12'b111111110011
;
      C0 <= 19'b0001110110100001101
;
      end
  7'd44:
     begin
      C1 <= 12'b111111110011
;
      C0 <= 19'b0001110000011010111
;
      end
  7'd45:
     begin
      C1 <= 12'b111111110011
;
      C0 <= 19'b0001101010001100111
;
      end
  7'd46:
     begin
      C1 <= 12'b111111110010
;
      C0 <= 19'b0001100011111000001
;
      end
  7'd47:
     begin
      C1 <= 12'b111111110010
;
      C0 <= 19'b0001011101011100100
;
      end
  7'd48:
     begin
      C1 <= 12'b111111110010
;
      C0 <= 19'b0001010110111010001
;
      end
  7'd49:
     begin
      C1 <= 12'b111111110010
;
      C0 <= 19'b0001010000010001011
;
      end
  7'd50:
     begin
      C1 <= 12'b111111110001
;
      C0 <= 19'b0001001001100010001
;
      end
  7'd51:
     begin
      C1 <= 12'b111111110001
;
      C0 <= 19'b0001000010101100100
;
      end
  7'd52:
     begin
      C1 <= 12'b111111110001
;
      C0 <= 19'b0000111011110000111
;
      end
  7'd53:
     begin
      C1 <= 12'b111111110001
;
      C0 <= 19'b0000110100101111010
;
      end
  7'd54:
     begin
      C1 <= 12'b111111110000
;
      C0 <= 19'b0000101101100111110
;
      end
  7'd55:
     begin
      C1 <= 12'b111111110000
;
      C0 <= 19'b0000100110011010100
;
      end
  7'd56:
     begin
      C1 <= 12'b111111110000
;
      C0 <= 19'b0000011111000111101
;
      end
  7'd57:
     begin
      C1 <= 12'b111111110000
;
      C0 <= 19'b0000010111101111011
;
      end
  7'd58:
     begin
      C1 <= 12'b111111101111
;
      C0 <= 19'b0000010000010001111
;
      end
  7'd59:
     begin
      C1 <= 12'b111111101111
;
      C0 <= 19'b0000001000101111010
;
      end
  7'd60:
     begin
      C1 <= 12'b111111101111
;
      C0 <= 19'b0000000001000111101
;
      end
  7'd61:
     begin
      C1 <= 12'b111111101111
;
      C0 <= 19'b0011111001011011010
;
      end
  7'd62:
     begin
      C1 <= 12'b111111101111
;
      C0 <= 19'b0011110001101010010
;
      end
  7'd63:
     begin
      C1 <= 12'b111111101110
;
      C0 <= 19'b0011101001110100101
;
      end
  7'd64:
     begin
      C1 <= 12'b111111101110
;
      C0 <= 19'b0011100001111010110
;
      end
  7'd65:
     begin
      C1 <= 12'b111111101110
;
      C0 <= 19'b0011011001111100101
;
      end
  7'd66:
     begin
      C1 <= 12'b111111101110
;
      C0 <= 19'b0011010001111010100
;
      end
  7'd67:
     begin
      C1 <= 12'b111111101101
;
      C0 <= 19'b0011001001110100100
;
      end
  7'd68:
     begin
      C1 <= 12'b111111101101
;
      C0 <= 19'b0011000001101010111
;
      end
  7'd69:
     begin
      C1 <= 12'b111111101101
;
      C0 <= 19'b0010111001011101110
;
      end
  7'd70:
     begin
      C1 <= 12'b111111101101
;
      C0 <= 19'b0010110001001101010
;
      end
  7'd71:
     begin
      C1 <= 12'b111111101101
;
      C0 <= 19'b0010101000111001101
;
      end
  7'd72:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0010100000100010111
;
      end
  7'd73:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0010011000001001011
;
      end
  7'd74:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0010001111101101010
;
      end
  7'd75:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0010000111001110101
;
      end
  7'd76:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0001111110101101110
;
      end
  7'd77:
     begin
      C1 <= 12'b111111101100
;
      C0 <= 19'b0001110110001010101
;
      end
  7'd78:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001101101100101101
;
      end
  7'd79:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001100100111111000
;
      end
  7'd80:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001011100010110101
;
      end
  7'd81:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001010011101101000
;
      end
  7'd82:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001001011000010000
;
      end
  7'd83:
     begin
      C1 <= 12'b111111101011
;
      C0 <= 19'b0001000010010110001
;
      end
  7'd84:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000111001101001011
;
      end
  7'd85:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000110000111100000
;
      end
  7'd86:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000101000001110001
;
      end
  7'd87:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000011111100000001
;
      end
  7'd88:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000010110110001111
;
      end
  7'd89:
     begin
      C1 <= 12'b111111101010
;
      C0 <= 19'b0000001110000011111
;
      end
  7'd90:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0000000101010110001
;
      end
  7'd91:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011100000100100110
;
      end
  7'd92:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011011010111010010
;
      end
  7'd93:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011010101001101110
;
      end
  7'd94:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011001111011111001
;
      end
  7'd95:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011001001101110100
;
      end
  7'd96:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0011000011111011111
;
      end
  7'd97:
     begin
      C1 <= 12'b111111101001
;
      C0 <= 19'b0010111110000111100
;
      end
  7'd98:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010111000010001001
;
      end
  7'd99:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010110010011001001
;
      end
  7'd100:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010101100011111011
;
      end
  7'd101:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010100110100011111
;
      end
  7'd102:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010100000100110111
;
      end
  7'd103:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010011010101000010
;
      end
  7'd104:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010010100101000001
;
      end
  7'd105:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010001110100110101
;
      end
  7'd106:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010001000100011110
;
      end
  7'd107:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0010000010011111100
;
      end
  7'd108:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0001111100011010001
;
      end
  7'd109:
     begin
      C1 <= 12'b111111101000
;
      C0 <= 19'b0001110110010011011
;
      end
  7'd110:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001110000001011101
;
      end
  7'd111:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001101010000010110
;
      end
  7'd112:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001100011111000110
;
      end
  7'd113:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001011101101101111
;
      end
  7'd114:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001010111100010001
;
      end
  7'd115:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001010001010101100
;
      end
  7'd116:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001001011001000001
;
      end
  7'd117:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0001000100111010000
;
      end
  7'd118:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000111110101011010
;
      end
  7'd119:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000111000011011110
;
      end
  7'd120:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000110010001011111
;
      end
  7'd121:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000101011111011100
;
      end
  7'd122:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000100101101010101
;
      end
  7'd123:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000011111011001011
;
      end
  7'd124:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000011001000111111
;
      end
  7'd125:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000010010110110001
;
      end
  7'd126:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000001100100100001
;
      end
  7'd127:
     begin
      C1 <= 12'b111111100111
;
      C0 <= 19'b0000000110010010001
;
      end

default:
begin
	C1 <= 12'b0;
	C0 <= 19'b0;
end
endcase
end
endmodule