`include "def.v"

module sqrt ( x_f,
			  polysel,
			  y_f);
input [30:0]x_f;
input polysel;
output [19:0]y_f;

wire [5 : 0]x_f_a;
wire [30:0]x_f_b;
wire [11:0]C1_12;
wire [19:0]C0_12;  						// coefficients of piecewise polynomial in interval [1,2) and [2,4)
wire [11:0]C1_24;
wire [19:0]C0_24;
wire [11:0]C1;
wire [19:0]C0;

assign x_f_a = x_f[30 : 25];
assign x_f_b = x_f[24 : 0] << 6;				// range reduction


sqrt_poly_1_2 sqrt_poly_1_2_0(	.x_f_a(x_f_a),
								.C1_o(C1_12),
								.C0_o(C0_12) );
								
sqrt_poly_2_4 sqrt_poly_2_4_0(	.x_f_a(x_f_a),
								.C1_o(C1_24),
								.C0_o(C0_24) );
								
assign C0 = (polysel == `TRUE)? C0_12:  C0_24;					// selects interval based on the the input provided
assign C1 = (polysel == `TRUE)? C1_12 : C0_24;

/*Multiplies the coefficients with the input and produces the output*/
myMultiplier_sqrt9	myMultiplier_sqrt9_0 (.x_f_b(x_f_b),
										  .C1(C1),
										  .C0(C0),
										  .y_f(y_f));					   


								

endmodule


/******************************* This module acts as the look up for the square root in interval [1,2) and outputs the required coefficients*****************************/

module sqrt_poly_1_2(	x_f_a,
						C1_o,
						C0_o );
input [5:0]x_f_a;
output  [11:0]C1_o;
output  [19:0]C0_o;

reg [11:0]C1;
reg [19:0]C0;

assign C1_o = C1;
assign C0_o = C0;

always @(*)
begin
case(x_f_a)

 6'd0:
     begin
      C1 <= 12'b000000100000
;
      C0 <= 20'b01000000001111111011
;
      end
 6'd1:
     begin
      C1 <= 12'b000000100000
;
      C0 <= 20'b01000001101110111101
;
      end
 6'd2:
     begin
      C1 <= 12'b000000011111
;
      C0 <= 20'b01000011001100110001
;
      end
 6'd3:
     begin
      C1 <= 12'b000000011111
;
      C0 <= 20'b01000100101001011011
;
      end
 6'd4:
     begin
      C1 <= 12'b000000011111
;
      C0 <= 20'b01000110000100111110
;
      end
 6'd5:
     begin
      C1 <= 12'b000000011111
;
      C0 <= 20'b01000111011111011011
;
      end
 6'd6:
     begin
      C1 <= 12'b000000011110
;
      C0 <= 20'b01001000111000110100
;
      end
 6'd7:
     begin
      C1 <= 12'b000000011110
;
      C0 <= 20'b01001010010001001011
;
      end
 6'd8:
     begin
      C1 <= 12'b000000011110
;
      C0 <= 20'b01001011101000100011
;
      end
 6'd9:
     begin
      C1 <= 12'b000000011110
;
      C0 <= 20'b01001100111110111100
;
      end
 6'd10:
     begin
      C1 <= 12'b000000011110
;
      C0 <= 20'b01001110010100011010
;
      end
 6'd11:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01001111101000111101
;
      end
 6'd12:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01010000111100100110
;
      end
 6'd13:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01010010001111011001
;
      end
 6'd14:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01010011100001010101
;
      end
 6'd15:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01010100110010011101
;
      end
 6'd16:
     begin
      C1 <= 12'b000000011101
;
      C0 <= 20'b01010110000010110010
;
      end
 6'd17:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01010111010010010100
;
      end
 6'd18:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01011000100001000110
;
      end
 6'd19:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01011001101111001000
;
      end
 6'd20:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01011010111100011100
;
      end
 6'd21:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01011100001001000011
;
      end
 6'd22:
     begin
      C1 <= 12'b000000011100
;
      C0 <= 20'b01011101010100111110
;
      end
 6'd23:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01011110100000001101
;
      end
 6'd24:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01011111101010110010
;
      end
 6'd25:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01100000110100101111
;
      end
 6'd26:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01100001111110000010
;
      end
 6'd27:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01100011000110101111
;
      end
 6'd28:
     begin
      C1 <= 12'b000000011011
;
      C0 <= 20'b01100100001110110101
;
      end
 6'd29:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01100101010110010101
;
      end
 6'd30:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01100110011101010000
;
      end
 6'd31:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01100111100011101000
;
      end
 6'd32:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01101000101001011100
;
      end
 6'd33:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01101001101110101101
;
      end
 6'd34:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01101010110011011100
;
      end
 6'd35:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01101011110111101010
;
      end
 6'd36:
     begin
      C1 <= 12'b000000011010
;
      C0 <= 20'b01101100111011011000
;
      end
 6'd37:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01101101111110100110
;
      end
 6'd38:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01101111000001010100
;
      end
 6'd39:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110000000011100100
;
      end
 6'd40:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110001000101010101
;
      end
 6'd41:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110010000110101010
;
      end
 6'd42:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110011000111100001
;
      end
 6'd43:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110100000111111011
;
      end
 6'd44:
     begin
      C1 <= 12'b000000011001
;
      C0 <= 20'b01110101000111111010
;
      end
 6'd45:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01110110000111011101
;
      end
 6'd46:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01110111000110100110
;
      end
 6'd47:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111000000101010011
;
      end
 6'd48:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111001000011100111
;
      end
 6'd49:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111010000001100010
;
      end
 6'd50:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111010111111000011
;
      end
 6'd51:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111011111100001011
;
      end
 6'd52:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111100111000111100
;
      end
 6'd53:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111101110101010100
;
      end
 6'd54:
     begin
      C1 <= 12'b000000011000
;
      C0 <= 20'b01111110110001010101
;
      end
 6'd55:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b01111111101100111111
;
      end
 6'd56:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000000101000010010
;
      end
 6'd57:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000001100011001111
;
      end
 6'd58:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000010011101110110
;
      end
 6'd59:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000011011000000111
;
      end
 6'd60:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000100010010000011
;
      end
 6'd61:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000101001011101011
;
      end
 6'd62:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000110000100111101
;
      end
 6'd63:
     begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b10000110111101111011
;
      end

default:
	  begin
	  C1 <= 12'b0;
	  C0 <= 20'b0;
	  end

endcase

end
endmodule


/******************************* This module acts as the look up for the square root in interval [2,4) and outputs the required coefficients*****************************/


module sqrt_poly_2_4(	x_f_a,
						C1_o,
						C0_o );
input [5:0]x_f_a;
output  [11:0]C1_o;
output  [19:0]C0_o;

reg [11:0]C1;
reg [19:0]C0;

assign C1_o = C1;
assign C0_o = C0;


always @(*)
begin
case(x_f_a)

6'd0:
      begin
      C1 <= 12'b000000010111
;
      C0 <= 20'b01011010110111001001
;
      end
6'd1:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01011100010000110010
;
      end
6'd2:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01011101101001011010
;
      end
6'd3:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01011111000001000011
;
      end
6'd4:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01100000010111101111
;
      end
6'd5:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01100001101101011111
;
      end
6'd6:
      begin
      C1 <= 12'b000000010110
;
      C0 <= 20'b01100011000010010101
;
      end
6'd7:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01100100010110010011
;
      end
6'd8:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01100101101001011010
;
      end
6'd9:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01100110111011101100
;
      end
6'd10:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01101000001101001010
;
      end
6'd11:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01101001011101110110
;
      end
6'd12:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01101010101101110001
;
      end
6'd13:
      begin
      C1 <= 12'b000000010101
;
      C0 <= 20'b01101011111100111100
;
      end
6'd14:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01101101001011011000
;
      end
6'd15:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01101110011001000110
;
      end
6'd16:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01101111100110001000
;
      end
6'd17:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01110000110010011111
;
      end
6'd18:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01110001111110001100
;
      end
6'd19:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01110011001001001111
;
      end
6'd20:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01110100010011101010
;
      end
6'd21:
      begin
      C1 <= 12'b000000010100
;
      C0 <= 20'b01110101011101011101
;
      end
6'd22:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01110110100110101010
;
      end
6'd23:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01110111101111010001
;
      end
6'd24:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111000110111010100
;
      end
6'd25:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111001111110110010
;
      end
6'd26:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111011000101101101
;
      end
6'd27:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111100001100000101
;
      end
6'd28:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111101010001111011
;
      end
6'd29:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111110010111010000
;
      end
6'd30:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b01111111011100000101
;
      end
6'd31:
      begin
      C1 <= 12'b000000010011
;
      C0 <= 20'b10000000100000011010
;
      end
6'd32:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000001100100010000
;
      end
6'd33:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000010100111100111
;
      end
6'd34:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000011101010100000
;
      end
6'd35:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000100101100111100
;
      end
6'd36:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000101101110111011
;
      end
6'd37:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000110110000011101
;
      end
6'd38:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10000111110001100100
;
      end
6'd39:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10001000110010010000
;
      end
6'd40:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10001001110010100000
;
      end
6'd41:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10001010110010010111
;
      end
6'd42:
      begin
      C1 <= 12'b000000010010
;
      C0 <= 20'b10001011110001110011
;
      end
6'd43:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10001100110000110110
;
      end
6'd44:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10001101101111100000
;
      end
6'd45:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10001110101101110010
;
      end
6'd46:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10001111101011101100
;
      end
6'd47:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010000101001001110
;
      end
6'd48:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010001100110011000
;
      end
6'd49:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010010100011001100
;
      end
6'd50:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010011011111101001
;
      end
6'd51:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010100011011110000
;
      end
6'd52:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010101010111100001
;
      end
6'd53:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010110010010111101
;
      end
6'd54:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10010111001110000011
;
      end
6'd55:
      begin
      C1 <= 12'b000000010001
;
      C0 <= 20'b10011000001000110101
;
      end
6'd56:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011001000011010010
;
      end
6'd57:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011001111101011011
;
      end
6'd58:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011010110111010000
;
      end
6'd59:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011011110000110010
;
      end
6'd60:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011100101010000000
;
      end
6'd61:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011101100010111100
;
      end
6'd62:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011110011011100100
;
      end
6'd63:
      begin
      C1 <= 12'b000000010000
;
      C0 <= 20'b10011111010011111011
;
	  end
default:
	  begin
	  C1 <= 12'b0;
	  C0 <= 20'b0;
	  end
endcase
end
endmodule

